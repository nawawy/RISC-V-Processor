module mem (
input bla
output blalala
....
)
