module regfile (
  input [31:0] writeData;
  input[4:0]  address;
  input writeEnable;
  output[31:0] readData;

  
  
  endmodule
)
