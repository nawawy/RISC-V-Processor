module imm_handler (
input bla
output blalala
....
)
