module pc(
  input[1:0] sel_pc;
   
  output[31:0] pc_out;
);


endmodule
