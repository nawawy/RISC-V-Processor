module mem (
  input [31:0] address, dataIN,
  output [31:0] memout,
  input clk
)
  
  
  
  endmodule;
)
