module imm_handler (
  input [31:0] instr;
  output [31:0] imm;
  input[2:0] ctrl;
  
....
)
