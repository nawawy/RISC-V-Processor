module alu(
  input [31:0] srca, srcb;
  input [5:0] alu_ctrl;
  
  output [31:0] alu_out;
  output branch_out;
);

endmodule
