module controlunit(
  input [31:0] instr;
  output [29:0] controls;

);



endmodule
