module immediatehandler (
input bla
output blalala
....
)
