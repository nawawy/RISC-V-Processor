module regfile (
input bla
output blalala
....
)
